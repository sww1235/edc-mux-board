library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mux8_1 is
  port (i : in std_logic_vector(7 downto 0);
        o : out std_logic;
        ctl : in std_logic_vector(2 downto 0));

end mux8_1;


architecture arch of mux8_1 is

begin

end arch;
