FPGA-I2C-Slave/I2C_slave.vhd