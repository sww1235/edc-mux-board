FPGA-I2C-Slave/I2C_slave_TB.vhd