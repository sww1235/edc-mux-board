
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


package fullmixer_pkg is
  type port_t is array (23 downto 0) of SIGNED(15 downto 0); -- port type for IO ports
  type ctl_port_array_t is array (23 downto 0) of port_t;
  type buffer_t is array (23 downto 0) of SIGNED(31 downto 0);
end package;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.fullmixer_pkg.all;

entity fullmixer is   -- 24x24 mixer matrix: 8 R IO, 8 L IO 8 mic IO
  port (i     : in  port_t;
        o     : out port_t;
        ctl   : in  ctl_port_array_t);



end fullmixer;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.fullmixer_pkg.all;

architecture Algorithmic of fullmixer is
  signal vo : buffer_t;

begin

  vo(0) <= ((i(0) * ctl(0)(0)) + (i(1) * ctl(0)(1)) + (i(2) * ctl(0)(2)) + (i(3) * ctl(0)(3))
          + (i(4) * ctl(0)(4)) + (i(5) * ctl(0)(5)) + (i(6) * ctl(0)(6)) + (i(7) * ctl(0)(7))
          + (i(8) * ctl(0)(8)) + (i(9) * ctl(0)(9)) + (i(10) * ctl(0)(10))
          + (i(11) * ctl(0)(11)) + (i(12) * ctl(0)(12)) + (i(13) * ctl(0)(13))
          + (i(14) * ctl(0)(14)) + (i(15) * ctl(0)(15)) + (i(16) * ctl(0)(16))
          + (i(17) * ctl(0)(17)) + (i(18) * ctl(0)(18)) + (i(19) * ctl(0)(19))
          + (i(20) * ctl(0)(20)) + (i(21) * ctl(0)(21)) + (i(22) * ctl(0)(22)) + (i(23) * ctl(0)(23)));

  vo(1) <= ((i(0) * ctl(1)(0)) + (i(1) * ctl(1)(1)) + (i(2) * ctl(1)(2)) + (i(3) * ctl(1)(3))
          + (i(4) * ctl(1)(4)) + (i(5) * ctl(1)(5)) + (i(6) * ctl(1)(6)) + (i(7) * ctl(1)(7))
          + (i(8) * ctl(1)(8)) + (i(9) * ctl(1)(9)) + (i(10) * ctl(1)(10))
          + (i(11) * ctl(1)(11)) + (i(12) * ctl(1)(12)) + (i(13) * ctl(1)(13))
          + (i(14) * ctl(1)(14)) + (i(15) * ctl(1)(15)) + (i(16) * ctl(1)(16))
          + (i(17) * ctl(1)(17)) + (i(18) * ctl(1)(18)) + (i(19) * ctl(1)(19))
          + (i(20) * ctl(1)(20)) + (i(21) * ctl(1)(21)) + (i(22) * ctl(1)(22)) + (i(23) * ctl(1)(23)));

  vo(2) <= ((i(0) * ctl(2)(0)) + (i(1) * ctl(2)(1)) + (i(2) * ctl(2)(2)) + (i(3) * ctl(2)(3))
          + (i(4) * ctl(2)(4)) + (i(5) * ctl(2)(5)) + (i(6) * ctl(2)(6)) + (i(7) * ctl(2)(7))
          + (i(8) * ctl(2)(8)) + (i(9) * ctl(2)(9)) + (i(10) * ctl(2)(10))
          + (i(11) * ctl(2)(11)) + (i(12) * ctl(2)(12)) + (i(13) * ctl(2)(13))
          + (i(14) * ctl(2)(14)) + (i(15) * ctl(2)(15)) + (i(16) * ctl(2)(16))
          + (i(17) * ctl(2)(17)) + (i(18) * ctl(2)(18)) + (i(19) * ctl(2)(19))
          + (i(20) * ctl(2)(20)) + (i(21) * ctl(2)(21)) + (i(22) * ctl(2)(22)) + (i(23) * ctl(2)(23)));

  vo(3) <= ((i(0) * ctl(3)(0)) + (i(1) * ctl(3)(1)) + (i(2) * ctl(3)(2)) + (i(3) * ctl(3)(3))
          + (i(4) * ctl(3)(4)) + (i(5) * ctl(3)(5)) + (i(6) * ctl(3)(6)) + (i(7) * ctl(3)(7))
          + (i(8) * ctl(3)(8)) + (i(9) * ctl(3)(9)) + (i(10) * ctl(3)(10))
          + (i(11) * ctl(3)(11)) + (i(12) * ctl(3)(12)) + (i(13) * ctl(3)(13))
          + (i(14) * ctl(3)(14)) + (i(15) * ctl(3)(15)) + (i(16) * ctl(3)(16))
          + (i(17) * ctl(3)(17)) + (i(18) * ctl(3)(18)) + (i(19) * ctl(3)(19))
          + (i(20) * ctl(3)(20)) + (i(21) * ctl(3)(21)) + (i(22) * ctl(3)(22)) + (i(23) * ctl(3)(23)));

  vo(4) <= ((i(0) * ctl(4)(0)) + (i(1) * ctl(4)(1)) + (i(2) * ctl(4)(2)) + (i(3) * ctl(4)(3))
          + (i(4) * ctl(4)(4)) + (i(5) * ctl(4)(5)) + (i(6) * ctl(4)(6)) + (i(7) * ctl(4)(7))
          + (i(8) * ctl(4)(8)) + (i(9) * ctl(4)(9)) + (i(10) * ctl(4)(10))
          + (i(11) * ctl(4)(11)) + (i(12) * ctl(4)(12)) + (i(13) * ctl(4)(13))
          + (i(14) * ctl(4)(14)) + (i(15) * ctl(4)(15)) + (i(16) * ctl(4)(16))
          + (i(17) * ctl(4)(17)) + (i(18) * ctl(4)(18)) + (i(19) * ctl(4)(19))
          + (i(20) * ctl(4)(20)) + (i(21) * ctl(4)(21)) + (i(22) * ctl(4)(22)) + (i(23) * ctl(4)(23)));

  vo(5) <= ((i(0) * ctl(5)(0)) + (i(1) * ctl(5)(1)) + (i(2) * ctl(5)(2)) + (i(3) * ctl(5)(3))
          + (i(4) * ctl(5)(4)) + (i(5) * ctl(5)(5)) + (i(6) * ctl(5)(6)) + (i(7) * ctl(5)(7))
          + (i(8) * ctl(5)(8)) + (i(9) * ctl(5)(9)) + (i(10) * ctl(5)(10))
          + (i(11) * ctl(5)(11)) + (i(12) * ctl(5)(12)) + (i(13) * ctl(5)(13))
          + (i(14) * ctl(5)(14)) + (i(15) * ctl(5)(15)) + (i(16) * ctl(5)(16))
          + (i(17) * ctl(5)(17)) + (i(18) * ctl(5)(18)) + (i(19) * ctl(5)(19))
          + (i(20) * ctl(5)(20)) + (i(21) * ctl(5)(21)) + (i(22) * ctl(5)(22)) + (i(23) * ctl(5)(23)));

  vo(6) <= ((i(0) * ctl(6)(0)) + (i(1) * ctl(6)(1)) + (i(2) * ctl(6)(2)) + (i(3) * ctl(6)(3))
          + (i(4) * ctl(6)(4)) + (i(5) * ctl(6)(5)) + (i(6) * ctl(6)(6)) + (i(7) * ctl(6)(7))
          + (i(8) * ctl(6)(8)) + (i(9) * ctl(6)(9)) + (i(10) * ctl(6)(10))
          + (i(11) * ctl(6)(11)) + (i(12) * ctl(6)(12)) + (i(13) * ctl(6)(13))
          + (i(14) * ctl(6)(14)) + (i(15) * ctl(6)(15)) + (i(16) * ctl(6)(16))
          + (i(17) * ctl(6)(17)) + (i(18) * ctl(6)(18)) + (i(19) * ctl(6)(19))
          + (i(20) * ctl(6)(20)) + (i(21) * ctl(6)(21)) + (i(22) * ctl(6)(22)) + (i(23) * ctl(6)(23)));

  vo(7) <= ((i(0) * ctl(7)(0)) + (i(1) * ctl(7)(1)) + (i(2) * ctl(7)(2)) + (i(3) * ctl(7)(3))
          + (i(4) * ctl(7)(4)) + (i(5) * ctl(7)(5)) + (i(6) * ctl(7)(6)) + (i(7) * ctl(7)(7))
          + (i(8) * ctl(7)(8)) + (i(9) * ctl(7)(9)) + (i(10) * ctl(7)(10))
          + (i(11) * ctl(7)(11)) + (i(12) * ctl(7)(12)) + (i(13) * ctl(7)(13))
          + (i(14) * ctl(7)(14)) + (i(15) * ctl(7)(15)) + (i(16) * ctl(7)(16))
          + (i(17) * ctl(7)(17)) + (i(18) * ctl(7)(18)) + (i(19) * ctl(7)(19))
          + (i(20) * ctl(7)(20)) + (i(21) * ctl(7)(21)) + (i(22) * ctl(7)(22)) + (i(23) * ctl(7)(23)));

  vo(8) <= ((i(0) * ctl(8)(0)) + (i(1) * ctl(8)(1)) + (i(2) * ctl(8)(2)) + (i(3) * ctl(8)(3))
          + (i(4) * ctl(8)(4)) + (i(5) * ctl(8)(5)) + (i(6) * ctl(8)(6)) + (i(7) * ctl(8)(7))
          + (i(8) * ctl(8)(8)) + (i(9) * ctl(8)(9)) + (i(10) * ctl(8)(10))
          + (i(11) * ctl(8)(11)) + (i(12) * ctl(8)(12)) + (i(13) * ctl(8)(13))
          + (i(14) * ctl(8)(14)) + (i(15) * ctl(8)(15)) + (i(16) * ctl(8)(16))
          + (i(17) * ctl(8)(17)) + (i(18) * ctl(8)(18)) + (i(19) * ctl(8)(19))
          + (i(20) * ctl(8)(20)) + (i(21) * ctl(8)(21)) + (i(22) * ctl(8)(22)) + (i(23) * ctl(8)(23)));

  vo(9) <= ((i(0) * ctl(9)(0)) + (i(1) * ctl(9)(1)) + (i(2) * ctl(9)(2)) + (i(3) * ctl(9)(3))
          + (i(4) * ctl(9)(4)) + (i(5) * ctl(9)(5)) + (i(6) * ctl(9)(6)) + (i(7) * ctl(9)(7))
          + (i(8) * ctl(9)(8)) + (i(9) * ctl(9)(9)) + (i(10) * ctl(9)(10))
          + (i(11) * ctl(9)(11)) + (i(12) * ctl(9)(12)) + (i(13) * ctl(9)(13))
          + (i(14) * ctl(9)(14)) + (i(15) * ctl(9)(15)) + (i(16) * ctl(9)(16))
          + (i(17) * ctl(9)(17)) + (i(18) * ctl(9)(18)) + (i(19) * ctl(9)(19))
          + (i(20) * ctl(9)(20)) + (i(21) * ctl(9)(21)) + (i(22) * ctl(9)(22)) + (i(23) * ctl(9)(23)));

  vo(10) <= ((i(0) * ctl(10)(0)) + (i(1) * ctl(10)(1)) + (i(2) * ctl(10)(2)) + (i(3) * ctl(10)(3))
          + (i(4) * ctl(10)(4)) + (i(5) * ctl(10)(5)) + (i(6) * ctl(10)(6)) + (i(7) * ctl(10)(7))
          + (i(8) * ctl(10)(8)) + (i(9) * ctl(10)(9)) + (i(10) * ctl(10)(10))
          + (i(11) * ctl(10)(11)) + (i(12) * ctl(10)(12)) + (i(13) * ctl(10)(13))
          + (i(14) * ctl(10)(14)) + (i(15) * ctl(10)(15)) + (i(16) * ctl(10)(16))
          + (i(17) * ctl(10)(17)) + (i(18) * ctl(10)(18)) + (i(19) * ctl(10)(19))
          + (i(20) * ctl(10)(20)) + (i(21) * ctl(10)(21)) + (i(22) * ctl(10)(22)) + (i(23) * ctl(10)(23)));

  vo(11) <= ((i(0) * ctl(11)(0)) + (i(1) * ctl(11)(1)) + (i(2) * ctl(11)(2)) + (i(3) * ctl(11)(3))
          + (i(4) * ctl(11)(4)) + (i(5) * ctl(11)(5)) + (i(6) * ctl(11)(6)) + (i(7) * ctl(11)(7))
          + (i(8) * ctl(11)(8)) + (i(9) * ctl(11)(9)) + (i(10) * ctl(11)(10))
          + (i(11) * ctl(11)(11)) + (i(12) * ctl(11)(12)) + (i(13) * ctl(11)(13))
          + (i(14) * ctl(11)(14)) + (i(15) * ctl(11)(15)) + (i(16) * ctl(11)(16))
          + (i(17) * ctl(11)(17)) + (i(18) * ctl(11)(18)) + (i(19) * ctl(11)(19))
          + (i(20) * ctl(11)(20)) + (i(21) * ctl(11)(21)) + (i(22) * ctl(11)(22)) + (i(23) * ctl(11)(23)));

  vo(12) <= ((i(0) * ctl(12)(0)) + (i(1) * ctl(12)(1)) + (i(2) * ctl(12)(2)) + (i(3) * ctl(12)(3))
          + (i(4) * ctl(12)(4)) + (i(5) * ctl(12)(5)) + (i(6) * ctl(12)(6)) + (i(7) * ctl(12)(7))
          + (i(8) * ctl(12)(8)) + (i(9) * ctl(12)(9)) + (i(10) * ctl(12)(10))
          + (i(11) * ctl(12)(11)) + (i(12) * ctl(12)(12)) + (i(13) * ctl(12)(13))
          + (i(14) * ctl(12)(14)) + (i(15) * ctl(12)(15)) + (i(16) * ctl(12)(16))
          + (i(17) * ctl(12)(17)) + (i(18) * ctl(12)(18)) + (i(19) * ctl(12)(19))
          + (i(20) * ctl(12)(20)) + (i(21) * ctl(12)(21)) + (i(22) * ctl(12)(22)) + (i(23) * ctl(12)(23)));

  vo(13) <= ((i(0) * ctl(13)(0)) + (i(1) * ctl(13)(1)) + (i(2) * ctl(13)(2)) + (i(3) * ctl(13)(3))
          + (i(4) * ctl(13)(4)) + (i(5) * ctl(13)(5)) + (i(6) * ctl(13)(6)) + (i(7) * ctl(13)(7))
          + (i(8) * ctl(13)(8)) + (i(9) * ctl(13)(9)) + (i(10) * ctl(13)(10))
          + (i(11) * ctl(13)(11)) + (i(12) * ctl(13)(12)) + (i(13) * ctl(13)(13))
          + (i(14) * ctl(13)(14)) + (i(15) * ctl(13)(15)) + (i(16) * ctl(13)(16))
          + (i(17) * ctl(13)(17)) + (i(18) * ctl(13)(18)) + (i(19) * ctl(13)(19))
          + (i(20) * ctl(13)(20)) + (i(21) * ctl(13)(21)) + (i(22) * ctl(13)(22)) + (i(23) * ctl(13)(23)));

  vo(14) <= ((i(0) * ctl(14)(0)) + (i(1) * ctl(14)(1)) + (i(2) * ctl(14)(2)) + (i(3) * ctl(14)(3))
          + (i(4) * ctl(14)(4)) + (i(5) * ctl(14)(5)) + (i(6) * ctl(14)(6)) + (i(7) * ctl(14)(7))
          + (i(8) * ctl(14)(8)) + (i(9) * ctl(14)(9)) + (i(10) * ctl(14)(10))
          + (i(11) * ctl(14)(11)) + (i(12) * ctl(14)(12)) + (i(13) * ctl(14)(13))
          + (i(14) * ctl(14)(14)) + (i(15) * ctl(14)(15)) + (i(16) * ctl(14)(16))
          + (i(17) * ctl(14)(17)) + (i(18) * ctl(14)(18)) + (i(19) * ctl(14)(19))
          + (i(20) * ctl(14)(20)) + (i(21) * ctl(14)(21)) + (i(22) * ctl(14)(22)) + (i(23) * ctl(14)(23)));

  vo(15) <= ((i(0) * ctl(15)(0)) + (i(1) * ctl(15)(1)) + (i(2) * ctl(15)(2)) + (i(3) * ctl(15)(3))
          + (i(4) * ctl(15)(4)) + (i(5) * ctl(15)(5)) + (i(6) * ctl(15)(6)) + (i(7) * ctl(15)(7))
          + (i(8) * ctl(15)(8)) + (i(9) * ctl(15)(9)) + (i(10) * ctl(15)(10))
          + (i(11) * ctl(15)(11)) + (i(12) * ctl(15)(12)) + (i(13) * ctl(15)(13))
          + (i(14) * ctl(15)(14)) + (i(15) * ctl(15)(15)) + (i(16) * ctl(15)(16))
          + (i(17) * ctl(15)(17)) + (i(18) * ctl(15)(18)) + (i(19) * ctl(15)(19))
          + (i(20) * ctl(15)(20)) + (i(21) * ctl(15)(21)) + (i(22) * ctl(15)(22)) + (i(23) * ctl(15)(23)));

  vo(16) <= ((i(0) * ctl(16)(0)) + (i(1) * ctl(16)(1)) + (i(2) * ctl(16)(2)) + (i(3) * ctl(16)(3))
          + (i(4) * ctl(16)(4)) + (i(5) * ctl(16)(5)) + (i(6) * ctl(16)(6)) + (i(7) * ctl(16)(7))
          + (i(8) * ctl(16)(8)) + (i(9) * ctl(16)(9)) + (i(10) * ctl(16)(10))
          + (i(11) * ctl(16)(11)) + (i(12) * ctl(16)(12)) + (i(13) * ctl(16)(13))
          + (i(14) * ctl(16)(14)) + (i(15) * ctl(16)(15)) + (i(16) * ctl(16)(16))
          + (i(17) * ctl(16)(17)) + (i(18) * ctl(16)(18)) + (i(19) * ctl(16)(19))
          + (i(20) * ctl(16)(20)) + (i(21) * ctl(16)(21)) + (i(22) * ctl(16)(22)) + (i(23) * ctl(16)(23)));

  vo(17) <= ((i(0) * ctl(17)(0)) + (i(1) * ctl(17)(1)) + (i(2) * ctl(17)(2)) + (i(3) * ctl(17)(3))
          + (i(4) * ctl(17)(4)) + (i(5) * ctl(17)(5)) + (i(6) * ctl(17)(6)) + (i(7) * ctl(17)(7))
          + (i(8) * ctl(17)(8)) + (i(9) * ctl(17)(9)) + (i(10) * ctl(17)(10))
          + (i(11) * ctl(17)(11)) + (i(12) * ctl(17)(12)) + (i(13) * ctl(17)(13))
          + (i(14) * ctl(17)(14)) + (i(15) * ctl(17)(15)) + (i(16) * ctl(17)(16))
          + (i(17) * ctl(17)(17)) + (i(18) * ctl(17)(18)) + (i(19) * ctl(17)(19))
          + (i(20) * ctl(17)(20)) + (i(21) * ctl(17)(21)) + (i(22) * ctl(17)(22)) + (i(23) * ctl(17)(23)));

  vo(18) <= ((i(0) * ctl(18)(0)) + (i(1) * ctl(18)(1)) + (i(2) * ctl(18)(2)) + (i(3) * ctl(18)(3))
          + (i(4) * ctl(18)(4)) + (i(5) * ctl(18)(5)) + (i(6) * ctl(18)(6)) + (i(7) * ctl(18)(7))
          + (i(8) * ctl(18)(8)) + (i(9) * ctl(18)(9)) + (i(10) * ctl(18)(10))
          + (i(11) * ctl(18)(11)) + (i(12) * ctl(18)(12)) + (i(13) * ctl(18)(13))
          + (i(14) * ctl(18)(14)) + (i(15) * ctl(18)(15)) + (i(16) * ctl(18)(16))
          + (i(17) * ctl(18)(17)) + (i(18) * ctl(18)(18)) + (i(19) * ctl(18)(19))
          + (i(20) * ctl(18)(20)) + (i(21) * ctl(18)(21)) + (i(22) * ctl(18)(22)) + (i(23) * ctl(18)(23)));


  vo(19) <= ((i(0) * ctl(19)(0)) + (i(1) * ctl(19)(1)) + (i(2) * ctl(19)(2)) + (i(3) * ctl(19)(3))
          + (i(4) * ctl(19)(4)) + (i(5) * ctl(19)(5)) + (i(6) * ctl(19)(6)) + (i(7) * ctl(19)(7))
          + (i(8) * ctl(19)(8)) + (i(9) * ctl(19)(9)) + (i(10) * ctl(19)(10))
          + (i(11) * ctl(19)(11)) + (i(12) * ctl(19)(12)) + (i(13) * ctl(19)(13))
          + (i(14) * ctl(19)(14)) + (i(15) * ctl(19)(15)) + (i(16) * ctl(19)(16))
          + (i(17) * ctl(19)(17)) + (i(18) * ctl(19)(18)) + (i(19) * ctl(19)(19))
          + (i(20) * ctl(19)(20)) + (i(21) * ctl(19)(21)) + (i(22) * ctl(19)(22)) + (i(23) * ctl(19)(23)));

  vo(20) <= ((i(0) * ctl(20)(0)) + (i(1) * ctl(20)(1)) + (i(2) * ctl(20)(2)) + (i(3) * ctl(20)(3))
          + (i(4) * ctl(20)(4)) + (i(5) * ctl(20)(5)) + (i(6) * ctl(20)(6)) + (i(7) * ctl(20)(7))
          + (i(8) * ctl(20)(8)) + (i(9) * ctl(20)(9)) + (i(10) * ctl(20)(10))
          + (i(11) * ctl(20)(11)) + (i(12) * ctl(20)(12)) + (i(13) * ctl(20)(13))
          + (i(14) * ctl(20)(14)) + (i(15) * ctl(20)(15)) + (i(16) * ctl(20)(16))
          + (i(17) * ctl(20)(17)) + (i(18) * ctl(20)(18)) + (i(19) * ctl(20)(19))
          + (i(20) * ctl(20)(20)) + (i(21) * ctl(20)(21)) + (i(22) * ctl(20)(22)) + (i(23) * ctl(20)(23)));

  vo(21) <= ((i(0) * ctl(21)(0)) + (i(1) * ctl(21)(1)) + (i(2) * ctl(21)(2)) + (i(3) * ctl(21)(3))
          + (i(4) * ctl(21)(4)) + (i(5) * ctl(21)(5)) + (i(6) * ctl(21)(6)) + (i(7) * ctl(21)(7))
          + (i(8) * ctl(21)(8)) + (i(9) * ctl(21)(9)) + (i(10) * ctl(21)(10))
          + (i(11) * ctl(21)(11)) + (i(12) * ctl(21)(12)) + (i(13) * ctl(21)(13))
          + (i(14) * ctl(21)(14)) + (i(15) * ctl(21)(15)) + (i(16) * ctl(21)(16))
          + (i(17) * ctl(21)(17)) + (i(18) * ctl(21)(18)) + (i(19) * ctl(21)(19))
          + (i(20) * ctl(21)(20)) + (i(21) * ctl(21)(21)) + (i(22) * ctl(21)(22)) + (i(23) * ctl(21)(23)));

  vo(22) <= ((i(0) * ctl(22)(0)) + (i(1) * ctl(22)(1)) + (i(2) * ctl(22)(2)) + (i(3) * ctl(22)(3))
          + (i(4) * ctl(22)(4)) + (i(5) * ctl(22)(5)) + (i(6) * ctl(22)(6)) + (i(7) * ctl(22)(7))
          + (i(8) * ctl(22)(8)) + (i(9) * ctl(22)(9)) + (i(10) * ctl(22)(10))
          + (i(11) * ctl(22)(11)) + (i(12) * ctl(22)(12)) + (i(13) * ctl(22)(13))
          + (i(14) * ctl(22)(14)) + (i(15) * ctl(22)(15)) + (i(16) * ctl(22)(16))
          + (i(17) * ctl(22)(17)) + (i(18) * ctl(22)(18)) + (i(19) * ctl(22)(19))
          + (i(20) * ctl(22)(20)) + (i(21) * ctl(22)(21)) + (i(22) * ctl(22)(22)) + (i(23) * ctl(22)(23)));

  vo(23) <= ((i(0) * ctl(22)(0)) + (i(1) * ctl(22)(1)) + (i(2) * ctl(22)(2)) + (i(3) * ctl(22)(3))
          + (i(4) * ctl(22)(4)) + (i(5) * ctl(22)(5)) + (i(6) * ctl(22)(6)) + (i(7) * ctl(22)(7))
          + (i(8) * ctl(22)(8)) + (i(9) * ctl(22)(9)) + (i(10) * ctl(22)(10))
          + (i(11) * ctl(22)(11)) + (i(12) * ctl(22)(12)) + (i(13) * ctl(22)(13))
          + (i(14) * ctl(22)(14)) + (i(15) * ctl(22)(15)) + (i(16) * ctl(22)(16))
          + (i(17) * ctl(22)(17)) + (i(18) * ctl(22)(18)) + (i(19) * ctl(22)(19))
          + (i(20) * ctl(22)(20)) + (i(21) * ctl(22)(21)) + (i(22) * ctl(22)(22)) + (i(23) * ctl(22)(23)));


  o(0) <= vo(0)(23 downto 8);
  o(1) <= vo(1)(23 downto 8);
  o(2) <= vo(2)(23 downto 8);
  o(3) <= vo(3)(23 downto 8);
  o(4) <= vo(4)(23 downto 8);
  o(5) <= vo(5)(23 downto 8);
  o(6) <= vo(6)(23 downto 8);
  o(7) <= vo(7)(23 downto 8);
  o(8) <= vo(8)(23 downto 8);
  o(9) <= vo(9)(23 downto 8);
  o(10) <= vo(10)(23 downto 8);
  o(11) <= vo(11)(23 downto 8);
  o(12) <= vo(12)(23 downto 8);
  o(13) <= vo(13)(23 downto 8);
  o(14) <= vo(14)(23 downto 8);
  o(15) <= vo(15)(23 downto 8);
  o(16) <= vo(16)(23 downto 8);
  o(17) <= vo(17)(23 downto 8);
  o(18) <= vo(18)(23 downto 8);
  o(19) <= vo(19)(23 downto 8);
  o(20) <= vo(20)(23 downto 8);
  o(21) <= vo(21)(23 downto 8);
  o(22) <= vo(22)(23 downto 8);
  o(23) <= vo(23)(23 downto 8);




end Algorithmic;
