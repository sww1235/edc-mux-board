FPGA-I2C-Slave/txt_util.vhd