
entity mixer is   -- 8x1 mixer
  port (i : in array(8 downto 0) of bit_vector(15 downto 0);
        ctl : in array(8 downto 0) of bit_vector(15 downto 0);
        o : out bit_vector(15 downto 0));


end mixer

architecture arch of mixer is


end arch
