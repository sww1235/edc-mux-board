FPGA-I2C-Slave/debounce.vhd